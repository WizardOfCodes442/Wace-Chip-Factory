library ieee;
use ieee.std_logic_1164.all;

entity half_sub is 
    port(a, c:in bit)