VHDL Code:
library ieee;
use ieee.std_logic_1164.all;

entity or1 is
    port(x, y)